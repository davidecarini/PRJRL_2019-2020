library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-----------------------------------------------------------------------
-- Unit�: Decoder_5_32
-- Descrizione: Decoder che trasforma una codifica binaria naturale in
-- una codifica one-hot.
-- Autore: Davide Carini
-----------------------------------------------------------------------
entity DECODER_5_32 is
generic( N_IN: INTEGER; N_OUT: INTEGER );
	port( 
		IN1:  IN  STD_LOGIC_VECTOR(N_IN-1 downto 0);
		OUT1: OUT STD_LOGIC_VECTOR(N_OUT -1 downto 0)
	);
end DECODER_5_32;

architecture RTL of DECODER_5_32 is

begin
	
  OUT1 <="00000000000000000000000000000001" when IN1="00000"else
         "00000000000000000000000000000010" when IN1="00001"else
         "00000000000000000000000000000100" when IN1="00010"else
         "00000000000000000000000000001000" when IN1="00011"else
			"00000000000000000000000000010000" when IN1="00100"else
			"00000000000000000000000000100000" when IN1="00101"else
			"00000000000000000000000001000000" when IN1="00110"else
			"00000000000000000000000010000000" when IN1="00111"else
			"00000000000000000000000100000000" when IN1="01000"else
			"00000000000000000000001000000000" when IN1="01001"else
			"00000000000000000000010000000000" when IN1="01010"else
			"00000000000000000000100000000000" when IN1="01011"else
			"00000000000000000001000000000000" when IN1="01100"else
			"00000000000000000010000000000000" when IN1="01101"else
			"00000000000000000100000000000000" when IN1="01110"else
			"00000000000000001000000000000000" when IN1="01111"else
			"00000000000000010000000000000000" when IN1="10000"else
			"00000000000000100000000000000000" when IN1="10001"else
			"00000000000001000000000000000000" when IN1="10010"else
			"00000000000010000000000000000000" when IN1="10011"else
			"00000000000100000000000000000000" when IN1="10100"else
			"00000000001000000000000000000000" when IN1="10101"else
			"00000000010000000000000000000000" when IN1="10110"else
			"00000000100000000000000000000000" when IN1="10111"else
			"00000001000000000000000000000000" when IN1="11000"else
			"00000010000000000000000000000000" when IN1="11001"else
			"00000100000000000000000000000000" when IN1="11010"else
			"00001000000000000000000000000000" when IN1="11011"else
			"00010000000000000000000000000000" when IN1="11100"else
			"00100000000000000000000000000000" when IN1="11101"else
			"01000000000000000000000000000000" when IN1="11110"else
			"10000000000000000000000000000000" when IN1="11111"else
			"--------------------------------" ;
end RTL;

